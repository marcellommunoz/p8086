library verilog;
use verilog.vl_types.all;
entity p8086 is
    port(
        clock           : in     vl_logic;
        reset           : in     vl_logic;
        wDEBUG          : in     vl_logic;
        entradaAX       : in     vl_logic_vector(15 downto 0);
        entradaBX       : in     vl_logic_vector(15 downto 0);
        entradaCX       : in     vl_logic_vector(15 downto 0);
        entradaDX       : in     vl_logic_vector(15 downto 0);
        entradaSP       : in     vl_logic_vector(15 downto 0);
        entradaBP       : in     vl_logic_vector(15 downto 0);
        entradaDI       : in     vl_logic_vector(15 downto 0);
        entradaSI       : in     vl_logic_vector(15 downto 0);
        entradaCS       : in     vl_logic_vector(15 downto 0);
        entradaDS       : in     vl_logic_vector(15 downto 0);
        entradaSS       : in     vl_logic_vector(15 downto 0);
        entradaES       : in     vl_logic_vector(15 downto 0);
        entradaIP       : in     vl_logic_vector(15 downto 0);
        entradaI1       : in     vl_logic_vector(15 downto 0);
        entradaI2       : in     vl_logic_vector(15 downto 0);
        entradaI3       : in     vl_logic_vector(15 downto 0);
        saidaAX         : out    vl_logic_vector(15 downto 0);
        saidaBX         : out    vl_logic_vector(15 downto 0);
        saidaCX         : out    vl_logic_vector(15 downto 0);
        saidaDX         : out    vl_logic_vector(15 downto 0);
        saidaSP         : out    vl_logic_vector(15 downto 0);
        saidaBP         : out    vl_logic_vector(15 downto 0);
        saidaDI         : out    vl_logic_vector(15 downto 0);
        saidaSI         : out    vl_logic_vector(15 downto 0);
        saidaCS         : out    vl_logic_vector(15 downto 0);
        saidaDS         : out    vl_logic_vector(15 downto 0);
        saidaSS         : out    vl_logic_vector(15 downto 0);
        saidaES         : out    vl_logic_vector(15 downto 0);
        saidaIP         : out    vl_logic_vector(15 downto 0);
        saidaI1         : out    vl_logic_vector(15 downto 0);
        saidaI2         : out    vl_logic_vector(15 downto 0);
        saidaI3         : out    vl_logic_vector(15 downto 0);
        SFROut          : out    vl_logic_vector(15 downto 0)
    );
end p8086;
