library verilog;
use verilog.vl_types.all;
entity p8086_vlg_vec_tst is
end p8086_vlg_vec_tst;
